/**
 * Copyright (C) 2025  AGH University of Science and Technology
 * 2025  AGH University of Science and Technology
 * MTM UEC2
 * Author: Dawid Bodzek
 *
 * Description:
 * Package with map related constants.
 */

package mapPkg;

    localparam LADDER_WIDTH = 32;
    localparam LADDER_HEIGHT = 32;
    localparam RAMP_OFFSET = 4;

    localparam LADDER_1_VSTART = 591;
    localparam LADDER_1_VSTOP = 716;
    localparam LADDER_1_HSTART = 796;
    localparam LADDER_1_HSTOP = 828;

    localparam LADDER_2_VSTART = 398;
    localparam LADDER_2_VSTOP = 567;
    localparam LADDER_2_HSTART = 388;
    localparam LADDER_2_HSTOP = 420;

    localparam LADDER_3_VSTART = 410;
    localparam LADDER_3_VSTOP = 555;
    localparam LADDER_3_HSTART = 196;
    localparam LADDER_3_HSTOP = 228;

    localparam LADDER_4_VSTART = 247;
    localparam LADDER_4_VSTOP = 372;
    localparam LADDER_4_HSTART = 796;
    localparam LADDER_4_HSTOP = 828;

    localparam LADDER_5_VSTART = 128;
    localparam LADDER_5_VSTOP = 271;
    localparam LADDER_5_HSTART = 544;
    localparam LADDER_5_HSTOP = 576;

endpackage