/**
 * Copyright (C) 2025  AGH University of Science and Technology
 * 2025  AGH University of Science and Technology
 * MTM UEC2
 * Author: Dawid Bodzek
 *
 * Description:
 * Package with ladder related constants.
 */

 package ladder_pkg;

    localparam LADDER_OFFSET = 16;
    localparam LADDER_WIDTH = 32;
    localparam LADDER_HEIGHT = 32;

    localparam LADDER_1_VSTART = 591;
    localparam LADDER_1_VSTOP = 716;
    localparam LADDER_1_HSTART = 796;

    localparam LADDER_2_VSTART = 398;
    localparam LADDER_2_VSTOP = 567;
    localparam LADDER_2_HSTART = 412;

    localparam LADDER_3_VSTART = 410;
    localparam LADDER_3_VSTOP = 555;
    localparam LADDER_3_HSTART = 220;

    localparam LADDER_4_VSTART = 247;
    localparam LADDER_4_VSTOP = 372;
    localparam LADDER_4_HSTART = 796;

    localparam LADDER_5_VSTART = 128;
    localparam LADDER_5_VSTOP = 271;
    localparam LADDER_5_HSTART = 544;

    localparam DECORATION_1_VSTART = 704;
    localparam DECORATION_1_VSTART_2 = 588;
    localparam DECORATION_1_HSTART = 320;

    localparam DECORATION_2_VSTART = 271;
    localparam DECORATION_2_VSTART_2 = 354;
    localparam DECORATION_2_HSTART = 576;

endpackage