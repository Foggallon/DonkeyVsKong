/**
 * Copyright (C) 2025  AGH University of Science and Technology
 * 2025  AGH University of Science and Technology
 * MTM UEC2
 * Author: Dawid Bodzek & Jakub Bukowski
 *
 * Description:
 * Package with kong character constants.
 */

package kong_pkg;

    localparam KONG_JUMP_HEIGHT = 58;
    localparam JUMP_TAKI_W_MIARE = 1_400_000;
    localparam MOVE_TAKI_NIE_MACQUEEN = 250_000;

    localparam KONG_ANIMATION_INITIAL_XPOS = 484;
    localparam KONG_ANIMATION_INITIAL_YPOS = 672;
    localparam KONG_PLATFORM_YPOS = 175;
    localparam KONG_PLATFORM_XPOS = 192;

    localparam CHARACTER_WIDTH = 64;
    localparam CHARACTER_HEIGHT = 64;

endpackage