/**
 * Copyright (C) 2025  AGH University of Science and Technology
 * MTM UEC2
 * Author: Dawid Bodzek
 *
 * Description:
 * Package with keyboard keys constants.
 */

package keyboard_pkg;

    localparam D = 'h3233;
    localparam A = 'h3143;
    localparam RELEASED = 'h4630;
    localparam SPACE = 'h3239;

endpackage