/**
 * San Jose State University
 * EE178 Lab #4
 * Author: prof. Eric Crabilla
 *
 * Modified by:
 * 2025  AGH University of Science and Technology
 * MTM UEC2
 * Piotr Kaczmarczyk
 *
 * Description:
 * Top level synthesizable module including the project top and all the FPGA-referred modules.
 */

module top_game_basys3 (
    input  wire clk,
    input  wire btnC,
    output wire Vsync,
    output wire Hsync,
    output wire [3:0] vgaRed,
    output wire [3:0] vgaGreen,
    output wire [3:0] vgaBlue,
    output wire JA1,

    inout wire PS2Clk,
    inout wire PS2Data
);

    timeunit 1ns;
    timeprecision 1ps;

    /**
     * Local variables and signals
     */

    wire clk40MHz;
    wire clk40MHz_mirror;
    wire clk100MHz;

    (* KEEP = "TRUE" *)
    (* ASYNC_REG = "TRUE" *)

    /**
     * Signals assignments
     */

    assign JA1 = clk40MHz_mirror;

    /**
     * FPGA submodules placement
     */

    clk_wiz_0 u_clk_wiz_0 (
        .clk,
        .clk100MHz,
        .clk40MHz,
        .locked()
    );

    ODDR pclk_oddr (
        .Q(clk40MHz_mirror),
        .C(clk40MHz),
        .CE(1'b1),
        .D1(1'b1),
        .D2(1'b0),
        .R(1'b0),
        .S(1'b0)
    );

    /**
     *  Project functional top module
     */

    top_game u_top_game (
        .clk40MHz,
        .clk100MHz,
        .ps2_clk(PS2Clk),
        .ps2_data(PS2Data),
        .rst(btnC),
        .r(vgaRed),
        .g(vgaGreen),
        .b(vgaBlue),
        .hs(Hsync),
        .vs(Vsync)
    );

endmodule