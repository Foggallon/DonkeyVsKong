/**
 * Copyright (C) 2025  AGH University of Science and Technology
 * 2025  AGH University of Science and Technology
 * MTM UEC2
 * Author: Dawid Bodzek
 *
 * Description:
 * Package with animation related constants.
 */

 package animation_pkg;

    localparam LADDER_VSTART = 271;
    localparam LADDER_HSTART = 480;
    localparam LADDER_HSTART_2 = 516;
    localparam PLATFORM_VSTART = 362;
    localparam PLATFORM_VSTART_2 = 539;

endpackage