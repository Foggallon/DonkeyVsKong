/**
 * Copyright (C) 2025  AGH University of Science and Technology
 * 2025  AGH University of Science and Technology
 * MTM UEC2
 * 
 * Author: Jakub Bukowski
 * Modified: Dawid Bodzek
 * 
 * Description:
 * The project top module.
 */

 module top_game (
   input  logic       clk65MHz,
   input  logic       rst,
   input  logic       ps2_clk,
   input  logic       ps2_data,
   output logic       vs,
   output logic       hs,
   output logic [3:0] r,
   output logic [3:0] g,
   output logic [3:0] b
);

   timeunit 1ns;
   timeprecision 1ps;

   /**
    * Interface definitions
    */

   vga_if draw_menu_if();
   vga_if vga_timing_if();
   vga_if draw_donkey_if();
   vga_if draw_ladder_if();
   vga_if platform_if();
   vga_if animation_ladder_if();
   vga_if animation_platform_if();
   vga_if draw_kong_if();
   vga_if draw_barrel_if();

   /**
    * Local variables and signals
    */

   logic animation;
   logic [3:0] counter, ctl;
   logic [11:0] rgb_pixel, rgb_pixel_menu, rgb_pixel_ladder, rgb_pixel_ramp, rgb_pixel_Aladder, rgb_pixel_Aramp, rgb_pixel_kong, rgb_pixel_barrel;
   logic [10:0] pixel_addr_ramp, pixel_addr_Aramp;
   logic [9:0] pixel_addr_ladder, pixel_addr_Aladder;
   logic [11:0] pixel_addr, pixel_addr_kong,  pixel_addr_barrel;
   logic [13:0] pixel_addr_menu;
   logic [10:0] xpos, ypos, xpos_kong, ypos_kong;

   logic [4:0] barrel;
   logic [4:0] barrel_v;
   logic done_1, done_2, done_3, done_4, done_5;
   logic done_ver_1, done_ver_2, done_ver_3, done_ver_4, done_ver_5;
   logic [9:0][10:0] xpos_barrel, ypos_barrel;
   logic [10:0] xpos_barrel_1, ypos_barrel_1, xpos_barrel_1_v, ypos_barrel_1_v;
   logic [10:0] xpos_barrel_2, ypos_barrel_2, xpos_barrel_2_v, ypos_barrel_2_v;
   logic [10:0] xpos_barrel_3, ypos_barrel_3, xpos_barrel_3_v, ypos_barrel_3_v;
   logic [10:0] xpos_barrel_4, ypos_barrel_4, xpos_barrel_4_v, ypos_barrel_4_v;
   logic [10:0] xpos_barrel_5, ypos_barrel_5, xpos_barrel_5_v, ypos_barrel_5_v;

   logic [15:0] keycode;
   logic [31:0] ascii_code;
   logic left, right, jump, rotate, start_game, up, down;

   /**
    * Signals assignments
    */

   assign xpos_barrel[0] = xpos_barrel_1;
   assign ypos_barrel[0] = ypos_barrel_1;
   assign xpos_barrel[1] = xpos_barrel_2;
   assign ypos_barrel[1] = ypos_barrel_2;
   assign xpos_barrel[2] = xpos_barrel_3;
   assign ypos_barrel[2] = ypos_barrel_3;
   assign xpos_barrel[3] = xpos_barrel_4;
   assign ypos_barrel[3] = ypos_barrel_4;
   assign xpos_barrel[4] = xpos_barrel_5;
   assign ypos_barrel[4] = ypos_barrel_5;
   assign xpos_barrel[5] = xpos_barrel_1_v;
   assign ypos_barrel[5] = ypos_barrel_1_v;
   assign xpos_barrel[6] = xpos_barrel_2_v;
   assign ypos_barrel[6] = ypos_barrel_2_v;
   assign xpos_barrel[7] = xpos_barrel_3_v;
   assign ypos_barrel[7] = ypos_barrel_3_v;
   assign xpos_barrel[8] = xpos_barrel_4_v;
   assign ypos_barrel[8] = ypos_barrel_4_v;
   assign xpos_barrel[9] = xpos_barrel_5_v;
   assign ypos_barrel[9] = ypos_barrel_5_v;

   assign vs = draw_donkey_if.vsync;
   assign hs = draw_donkey_if.hsync;
   assign {r,g,b} = draw_donkey_if.rgb;
   
   /**
    * Submodules instances
    */

   ps2_receiver u_ps2_receiver (
      .clk(clk65MHz),
      .kclk(ps2_clk),
      .kdata(ps2_data),
      .keycode(keycode),
      .oflag()
   );       

   bin2ascii u_bin2ascii (
      .I(keycode),
      .O(ascii_code)
  );

  key_decoder u_key_decoder (
      .clk(clk65MHz),
      .rst,
      .left,
      .right,
      .jump,
      .start_game(start_game),
      .up,
      .down,
      .keyCode(ascii_code),
      .rotate
   );

   vga_timing u_vga_timing (
      .clk(clk65MHz),
      .rst,
      
      .out(vga_timing_if)
  );

  image_rom  #(
      .BITS(14),
      .PIXELS(12292),
      .ROM_FILE("../../rtl/MainMenu/DonkeyVsKong_small.dat")
   ) u_image_Rom_menu (
      .clk(clk65MHz),
      .address(pixel_addr_menu),
      .rgb(rgb_pixel_menu)
   );

   draw_menu u_draw_menu (
      .clk(clk65MHz),
      .rst,
      .start_game,
      .pixel_addr(pixel_addr_menu),
      .rgb_pixel(rgb_pixel_menu),

      .in(vga_timing_if),
      .out(draw_menu_if)
   );

   animation_ladder u_animation_ladder (
        .clk(clk65MHz),
        .rst,
        .pixel_addr(pixel_addr_Aladder),
        .rgb_pixel(rgb_pixel_Aladder),
        .start_game,
        .animation,
        .counter(counter),
        .in(animation_platform_if),
        .out(animation_ladder_if)
   );

   image_rom  #(
        .BITS(10),
        .PIXELS(1028),
        .ROM_FILE("../../rtl/LevelElements/drabinka.dat")
    ) u_image_rom_Aladder (
      .clk(clk65MHz),
      .address(pixel_addr_Aladder),
      .rgb(rgb_pixel_Aladder)
   );

   animation_platform u_animation_platform (
        .clk(clk65MHz),
        .rst,
        .pixel_addr(pixel_addr_Aramp),
        .rgb_pixel(rgb_pixel_Aramp),
        .start_game,
        .ctl(ctl),
        .in(platform_if),
        .out(animation_platform_if)
    );

    image_rom  #(
        .BITS(11),
        .PIXELS(2052),
        .ROM_FILE("../../rtl/LevelElements/platforma.dat")
   ) u_image_rom_Aplatform (
      .clk(clk65MHz),
      .address(pixel_addr_Aramp),
      .rgb(rgb_pixel_Aramp)
   );

   start_animation u_start_animation (
      .clk(clk65MHz),
      .rst,
      .start_game,
      .animation(animation),
      .counter,
      .ctl,
      .xpos(xpos_kong),
      .ypos(ypos_kong)
   );

   draw_character #(
      .CHARACTER_HEIGHT(64),
      .CHARACTER_WIDTH(64)
   ) u_draw_character_kong (
      .clk(clk65MHz),
      .rst,
      .rotate('0),
      .start_game,
      .pixel_addr(pixel_addr_kong),
      .rgb_pixel(rgb_pixel_kong),
      .xpos(xpos_kong),
      .ypos(ypos_kong),
      .en(animation),

      .in(animation_ladder_if),
      .out(draw_kong_if)
   );
   
   image_rom  #(
      .BITS(12),
      .PIXELS(4096),
      .ROM_FILE("../../rtl/Kong/Kong.dat")
   
   ) u_image_rom_kong (
      .clk(clk65MHz),
      .address(pixel_addr_kong),
      .rgb(rgb_pixel_kong)
   );

   draw_ladder u_draw_ladder (
      .clk(clk65MHz),
      .rst,
      .start_game,
      .animation,
      .pixel_addr(pixel_addr_ladder),
      .rgb_pixel(rgb_pixel_ladder),

      .in(draw_menu_if),
      .out(draw_ladder_if)
   );

   image_rom  #(
        .BITS(10),
        .PIXELS(1028),
        .ROM_FILE("../../rtl/LevelElements/drabinka.dat")
   ) u_image_rom_ladder (
      .clk(clk65MHz),
      
      .address(pixel_addr_ladder),
      .rgb(rgb_pixel_ladder)
   );

   incline_platform u_incline_platform (
      .clk(clk65MHz),
      .rst,
      .pixel_addr(pixel_addr_ramp),
      .rgb_pixel(rgb_pixel_ramp),
      .start_game,
      .ctl,

      .in(draw_ladder_if),
      .out(platform_if)
   );

   image_rom  #(
      .BITS(11),
      .PIXELS(2052),
      .ROM_FILE("../../rtl/LevelElements/platforma.dat")
   ) u_image_rom_platform (
      .clk(clk65MHz),
      .address(pixel_addr_ramp),
      .rgb(rgb_pixel_ramp)
   );

   draw_character #(
      .CHARACTER_HEIGHT(64),
      .CHARACTER_WIDTH(48)
   ) u_draw_character_donkey (
      .clk(clk65MHz),
      .rst,
      .rotate,
      .start_game,
      .pixel_addr,
      .rgb_pixel,
      .xpos(xpos),
      .ypos(ypos),
      .en(!animation),

      .in(draw_barrel_if),
      .out(draw_donkey_if)
   );
   
   image_rom  #(
      .BITS(12),
      .PIXELS(4096),
      .ROM_FILE("../../rtl/Donkey/Donkey_v1.dat")
   
   ) u_image_rom_donkey (
      .clk(clk65MHz),
      
      .address(pixel_addr),
      .rgb(rgb_pixel)
   );

   donkey_movement u_donkey_movement (
      .clk(clk65MHz),
      .rst(rst),
      .xpos(xpos),
      .ypos(ypos),
      
      .start_game,
      .animation,
      .left,
      .right,
      .jump,
      .down,
      .up
   );

   hor_barrel u_ver_barrel_1 (
      .clk(clk65MHz),
      .rst(rst),
      .barrel(barrel[0]),
      .done(done_1),
      .xpos(xpos_barrel_1),
      .ypos(ypos_barrel_1)
   );

   hor_barrel u_ver_barrel_2 (
      .clk(clk65MHz),
      .rst(rst),
      .barrel(barrel[1]),
      .done(done_2),
      .xpos(xpos_barrel_2),
      .ypos(ypos_barrel_2)
   );

   hor_barrel u_ver_barrel_3 (
      .clk(clk65MHz),
      .rst(rst),
      .barrel(barrel[2]),
      .done(done_3),
      .xpos(xpos_barrel_3),
      .ypos(ypos_barrel_3)
   );

   hor_barrel u_ver_barrel_4 (
      .clk(clk65MHz),
      .rst(rst),
      .barrel(barrel[3]),
      .done(done_4),
      .xpos(xpos_barrel_4),
      .ypos(ypos_barrel_4)
   );

   hor_barrel u_ver_barrel_5 (
      .clk(clk65MHz),
      .rst(rst),
      .barrel(barrel[4]),
      .done(done_5),
      .xpos(xpos_barrel_5),
      .ypos(ypos_barrel_5)
   );

   ver_barrel u_ver_barrel_1_v (
      .clk(clk65MHz),
      .rst(rst),
      .xpos_kong(xpos_kong),
      .barrel(barrel_v[0]),
      .done(done_ver_1),
      .xpos(xpos_barrel_1_v),
      .ypos(ypos_barrel_1_v)
   );

   ver_barrel u_ver_barrel_2_v (
      .clk(clk65MHz),
      .rst(rst),
      .xpos_kong(xpos_kong),
      .barrel(barrel_v[1]),
      .done(done_ver_2),
      .xpos(xpos_barrel_2_v),
      .ypos(ypos_barrel_2_v)
   );

   ver_barrel u_ver_barrel_3_v (
      .clk(clk65MHz),
      .rst(rst),
      .xpos_kong(xpos_kong),
      .barrel(barrel_v[2]),
      .done(done_ver_3),
      .xpos(xpos_barrel_3_v),
      .ypos(ypos_barrel_3_v)
   );

   ver_barrel u_ver_barrel_4_v (
      .clk(clk65MHz),
      .rst(rst),
      .xpos_kong(xpos_kong),
      .barrel(barrel_v[3]),
      .done(done_ver_4),
      .xpos(xpos_barrel_4_v),
      .ypos(ypos_barrel_4_v)
   );

   ver_barrel u_ver_barrel_5_v (
      .clk(clk65MHz),
      .rst(rst),
      .xpos_kong(xpos_kong),
      .barrel(barrel_v[4]),
      .done(done_ver_5),
      .xpos(xpos_barrel_5_v),
      .ypos(ypos_barrel_5_v)
   );

   barrel_ctl #(.BARRELS(5), .DELAY_TIME(162_500_000)) u_barrel_ctl_hor (
      .clk(clk65MHz),
      .rst(rst),
      .start_game,
      .animation,
      .key(down),
      .done({done_5, done_4, done_3, done_2, done_1}),
      .barrel(barrel)
   );
   
   barrel_ctl #(.BARRELS(5), .DELAY_TIME(20_500_000)) u_barrel_ctl_ver (
      .clk(clk65MHz),
      .rst(rst),
      .start_game,
      .animation,
      .key(up),
      .done({done_ver_5, done_ver_4, done_ver_3, done_ver_2, done_ver_1}),
      .barrel(barrel_v)
   );

   draw_barrel #(.BARRELS(10)) u_draw_barrel (
      .clk(clk65MHz),
      .rst(rst),
      .start_game,
      .animation,
      .barrel({barrel_v, barrel}),
      .xpos(xpos_barrel),
      .ypos(ypos_barrel),
      .rgb_pixel(rgb_pixel_barrel),
      .pixel_addr(pixel_addr_barrel),

      .in(draw_kong_if),
      .out(draw_barrel_if)
   );

   image_rom  #(
      .BITS(12),
      .PIXELS(4096),
      .ROM_FILE("../../rtl/Donkey/Donkey_v1.dat")
   ) u_image_rom_barrel (
      .clk(clk65MHz),
      
      .address(pixel_addr_barrel),
      .rgb(rgb_pixel_barrel)
   );

endmodule