/**
 * Copyright (C) 2025  AGH University of Science and Technology
 * 2025  AGH University of Science and Technology
 * MTM UEC2
 * Author: Dawid Bodzek
 *
 * Description:
 * Package with barrel related constants.
 */

 package barrel_pkg;

    localparam BARREL_WIDTH = 32;
    localparam BARREL_HEIGHT = 32;
    localparam HOR_BARREL_INITIAL_YPOS = 208;
    localparam HIT_OFFSET = 4;
endpackage