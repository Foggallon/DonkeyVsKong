/**
 * Copyright (C) 2025  AGH University of Science and Technology
 * 2025  AGH University of Science and Technology
 * MTM UEC2
 * Author: Dawid Bodzek
 *
 * Description:
 * Package with donkey character constants.
 */

 package donkey_pkg;

    localparam DONKEY_JUMP_HEIGHT = 58;
    localparam JUMP_TAKI_W_MIARE = 1_400_000;
    localparam MOVE_TAKI_NIE_MACQUEEN = 250_000;

    localparam CHARACTER_HEIGHT = 64;
    localparam CHARACTER_WIDTH = 48;

    localparam DONKEY_INITIAL_XPOS = 128;
    localparam DONKEY_INITIAL_YPOS = 672;

endpackage